;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NGVD29
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements: 1166
652614.7178514417 4172927.2391306665  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "1_0"
652508.9283354593 4174610.913022432  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "1_1"
652822.3937414596 4175225.666186792  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "2_0"
652741.8734235434 4176148.585482046  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "2_1"
651463.2567447106 4175569.0074347947  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "3_0"
650572.1152749114 4176545.514108853  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "3_1"
650375.4934866645 4177467.8752769195  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "4_0"
650423.6788652857 4178227.182548184  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "4_1"
649544.2067746622 4180007.101882065  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "5_0"
649565.0228215281 4182305.052083309  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "5_1"
649531.827697602 4183060.253504173  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "6_0"
649281.2914525591 4183520.420989356  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "6_1"
648763.8612226166 4184776.937447396  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "7_0"
647656.4297185474 4185651.1804112205  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "7_1"
647397.3331177037 4185934.563526705  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "8_0"
648035.2836630072 4186190.02876331  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "8_1"
648246.3844216425 4187398.813136544  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "8_2"
648622.9734168162 4188933.923218364  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "9_0"
647700.8769792581 4190094.6571607674  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "9_1"
647585.3581625737 4190829.478914215  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "10_0"
647964.8535663108 4191302.2922414215  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "10_1"
647063.3913093798 4192798.1722151004  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "11_0"
646738.3811113861 4193826.493062018  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "11_1"
647100.7724014329 4194977.972240924  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "11_2"
647235.0011897258 4195628.583649331  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "12_0"
647323.2860568011 4197268.184213412  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "12_1"
647333.1467826745 4198957.44905271  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "13_0"
647021.09977915 4199766.549195513  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "14_0"
645786.190000817 4200284.775903742  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "15_0"
645966.6779999408 4201159.893432688  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "16_0"
646219.5219098359 4201426.458397796  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "16_1"
654339.4347903513 4171053.517097676  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "17_0"
653519.4837622403 4171454.228997129  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "17_1"
652699.6780225058 4171765.1027778825  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "17_2"
646034.0497289186 4201926.173677682  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "18_0"
645425.7151273586 4202115.77033329  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "18_1"
644985.7150489242 4202355.868746084  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "19_0"
644484.5130499462 4202604.326661308  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "19_1"
643713.6662048836 4203064.750156754  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "20_0"
642707.6742371497 4204210.731871361  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "21_0"
641783.1241133863 4205091.319808378  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "22_0"
641054.8322265873 4205642.276378543  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "22_1"
640116.1437944212 4206125.918347927  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "23_0"
639037.0220528527 4206574.849410551  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "24_0"
637997.2180230065 4206255.643113023  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "24_1"
637081.4248179944 4206612.490617054  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "25_0"
636541.1876787738 4207064.424014691  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "26_0"
636654.5552536811 4207423.611727671  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "26_1"
636875.1873247384 4207805.767230784  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "26_2"
635350.4745162827 4207356.338455758  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "27_0"
635674.0652994235 4207173.881105242  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "27_1"
635890.994157577 4207105.324961082  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "27_2"
636551.5141361423 4207953.036781178  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "28_0"
636141.2873738301 4208180.302101987  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "28_1"
635692.3887301612 4208357.545816318  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "28_2"
635519.9055204288 4208815.963231117  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "28_3"
635330.6522597591 4208099.76057296  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "29_0"
635201.9737194309 4207794.117685258  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "29_1"
635208.1652324264 4207480.319186943  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "29_2"
635824.2279465451 4207892.709324654  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "30_0"
635334.1207860553 4208729.886560926  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "31_0"
635112.5527831968 4209017.844299727  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "31_1"
634858.5556575002 4209392.497681738  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "31_2"
634519.1412973078 4209810.1655681105  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "31_3"
634403.7925257619 4209894.357213727  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "31_4"
633873.6211497841 4209717.824757041  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "32_0"
633500.4753748692 4209561.976678076  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "32_1"
632876.9697057205 4209972.18048305  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "32_2"
632442.7840635681 4210799.4817781085  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "33_0"
633285.8530504587 4210744.429387682  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "34_0"
632088.8742879326 4210861.580402396  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "35_0"
631778.96329538 4211106.041210271  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "35_1"
631385.1608874588 4211398.130439815  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "35_2"
631385.0422105627 4211677.233914774  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "35_3"
632593.2200627903 4211176.012888301  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "36_0"
632202.0512073531 4211454.343768115  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "36_1"
631993.2162240259 4211590.234754035  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "36_2"
631732.8605704183 4211860.7404659325  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "36_3"
631475.7299605195 4212071.807919479  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "36_4"
631472.3118061582 4212335.500938396  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "37_0"
630300.8748127669 4213017.163432803  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "37_1"
629685.0720415934 4213090.132817923  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "38_0"
629092.3120439798 4213160.263929328  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "38_1"
629078.7124956485 4213264.585295115  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "39_0"
628767.9415014661 4214634.935925243  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "40_0"
627812.9637436179 4213433.571722245  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "40_1"
628360.9648005284 4213193.388370545  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "41_0"
627799.6918708327 4213301.775114943  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "41_1"
626715.3125678551 4213653.73223194  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "42_0"
626825.7505163455 4213517.189673375  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "42_1"
626971.5182598662 4214671.365968964  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "42_2"
626517.0973087271 4215095.777965141  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "42_3"
626171.5160025129 4215543.254769776  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "42_4"
625775.7881344506 4215581.349289572  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "42_5"
625592.6591972457 4215838.780833752  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "43_0"
625636.6831789651 4216057.433030982  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "43_1"
625546.6405388041 4216443.278536714  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "44_0"
625363.8723625138 4217064.959026141  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "44_1"
625012.809920838 4217947.962649568  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "45_0"
624120.540799048 4218541.9983843705  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "45_1"
623354.0699693925 4218403.417849549  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "45_2"
622632.5401336574 4218787.022392843  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "45_3"
621811.2841889139 4217753.1418655915  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "45_4"
621361.220112684 4217500.240569754  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "46_0"
620888.4488036622 4217557.729687997  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "46_1"
620778.6565194229 4217247.233344266  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "46_2"
620778.6907216017 4216790.752048137  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "46_3"
620068.5017751172 4216135.677172261  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "46_4"
619480.9657340612 4216815.762449477  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "46_5"
619078.0452793605 4216911.07105481  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "46_6"
618884.1138476129 4217267.919545561  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "47_0"
618365.2015754777 4217297.731026506  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "47_1"
618075.1562609341 4217539.85145266  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "47_2"
617525.6530307748 4217710.285106714  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "47_3"
617006.0945918146 4216816.749289133  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "47_4"
616728.4228590499 4216762.273653913  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "47_5"
616430.814660026 4216644.658568676  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "47_6"
616193.5826177818 4216425.548048779  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "47_7"
616063.3558039457 4215684.9773234455  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "48_0"
616303.0309844827 4214745.106468371  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "48_1"
616284.7785602189 4214047.451553196  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "48_2"
614856.9309143114 4211089.157934559  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "49_0"
614007.652716993 4210171.271153342  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "49_1"
612403.2846640839 4209825.450978849  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "49_2"
611749.7603428664 4209709.297996088  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "49_3"
611621.7313268366 4209387.057954427  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "50_0"
609851.2989826737 4208742.540620985  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "50_1"
608835.6093210281 4209884.051282795  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "50_2"
608467.1418814643 4208733.846056663  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "51_0"
607763.639618161 4208373.831586166  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "51_1"
606606.4186983466 4208163.851360205  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "51_2"
605805.1267064564 4208896.47513682  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "51_3"
604988.5757998166 4208292.437865138  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "52_0"
604414.4645473409 4208347.405659039  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "52_1"
603946.5995082532 4209299.503574458  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "52_2"
603655.6071851981 4209660.46743191  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "52_3"
603324.9423712506 4209737.49223491  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "52_4"
603096.6526515429 4209890.082948687  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "52_5"
602523.7731173887 4210047.201161128  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_0"
602451.7517905527 4210250.455965163  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_1"
602288.7245001845 4210755.598632445  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_2"
602211.7564094145 4211053.610448057  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_3"
602164.6637928758 4211437.706040749  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_4"
602119.7778607586 4211742.873917756  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_5"
601993.4723119023 4212059.5807839595  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_6"
601990.9134244871 4212324.015319652  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_7"
601868.3859638646 4212550.516462428  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_8"
601833.0205114698 4212783.483337573  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "53_9"
646937.8381330459 4185892.7927735206  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "54_0"
646694.330867206 4185980.7560972613  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "54_1"
646643.7824279584 4186242.5411841287  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "54_2"
646818.7999934455 4186906.48532669  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "55_0"
646548.1575074961 4187276.0239843465  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "55_1"
646141.2301657741 4187070.2039506924  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "56_0"
645625.0797538795 4187239.130133253  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "56_1"
645374.8887557762 4187056.3878553538  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "57_0"
644678.819488807 4186877.158089837  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "57_1"
643939.1714584498 4186869.7720620125  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "58_0"
643287.045457815 4187165.1031422312  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "58_1"
643002.4764438212 4187363.4325330663  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "59_0"
642854.7376746334 4187140.809724125  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "59_1"
642598.035322276 4186660.487820532  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "60_0"
642437.992004464 4186377.730306525  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "60_1"
642016.6694409396 4185987.5091518327  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "60_2"
641515.1469174129 4185762.2708318117  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "61_0"
641224.4894858535 4185748.740583315  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "61_1"
640450.3222122159 4185530.7315101144  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "61_2"
640087.6540549084 4185799.5407181885  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "62_0"
639826.3143737331 4185988.9528127746  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "62_1"
639474.2818268305 4186170.626129978  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "62_2"
639336.8704274953 4185751.374429547  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "63_0"
639244.7974410157 4185497.4782129456  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "63_1"
639189.9253467575 4185224.0706555457  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "63_2"
639582.9903173889 4185651.9596389397  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "65_0"
639373.7917661609 4185947.092739678  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "65_1"
639423.6833469948 4185295.1773140384  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "66_0"
639259.5221554051 4185260.970633459  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "66_1"
639087.7752779205 4184981.1987560396  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "67_0"
638554.0294231656 4184151.8348933905  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "68_0"
638069.4186927608 4184217.5208286257  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "68_1"
638429.0453655269 4185046.490250335  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "69_0"
638054.1920484812 4184652.012388286  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "69_1"
637929.9940507486 4184625.7954040137  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "70_0"
637428.2848508954 4184873.2045919616  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "70_1"
636491.1761195434 4185454.499272559  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "71_0"
635884.4449167945 4184802.1393525978  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "71_1"
635178.4469824474 4185059.7707308363  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "72_0"
635063.8479694315 4184654.7381303087  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "72_1"
634973.4998721435 4184227.6296727965  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "73_0"
634572.5994903009 4183733.698621285  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "73_1"
634377.8473394773 4183518.4759107917  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "73_2"
633981.4067408236 4183076.6305899126  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "74_0"
633812.7577762684 4182742.526895528  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "74_1"
633079.4137154359 4182774.242766127  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "75_0"
632386.8073160099 4182769.634358488  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "75_1"
631811.7553594916 4183191.465963721  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "76_0"
631343.9402646346 4183665.1552534667  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "77_0"
630633.6657147555 4184008.09064878  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "77_1"
630124.0966504012 4184583.337684652  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "77_2"
629319.559581462 4185080.908353555  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "78_0"
628840.575746778 4185609.054718785  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "79_0"
628228.445779227 4186007.7100935974  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "80_0"
627423.013035264 4186402.4153376142  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "80_1"
627308.0277616375 4186602.721113504  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "81_0"
627541.9482293101 4187836.3286579642  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "82_0"
615682.4277215751 4212911.243595765  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "83_0"
615193.3915731206 4212529.25441579  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "83_1"
614948.1357014917 4212045.5780361695  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "83_2"
626956.483912094 4189824.5720677786  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "85_0"
626193.5846408063 4190937.482642918  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "86_0"
625603.3511694361 4191953.381675128  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "86_1"
625604.0246774505 4191989.324563052  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "88_0"
625123.7928637639 4192413.64304921  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "88_1"
625506.1848645561 4194056.0073785298  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "89_0"
625503.5421683704 4194390.986399873  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "90_0"
626142.2872272825 4195635.054212464  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "91_0"
625683.7702274414 4196105.7048  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "92_0"
626335.7184695086 4197325.990044627  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "94_0"
626618.3383862565 4197759.761262759  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "94_1"
626825.5314435746 4198829.212785309  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "95_0"
626548.1090363426 4199791.073976104  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "96_0"
626336.2774819357 4200522.0043511465  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "97_0"
626695.3372005516 4200422.026525206  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "98_0"
626555.5541922717 4200581.745482544  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "99_0"
626702.8179155738 4201230.459615269  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "100_0"
626428.8156815215 4201628.334261918  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "100_1"
625914.4713866932 4200723.637421671  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "101_0"
626176.0230869557 4201323.499414929  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "101_1"
625775.6960542941 4201619.919383359  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "102_0"
626320.5373437743 4202011.7762705535  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "103_0"
625315.8589383338 4201869.544247121  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "104_0"
625811.8421550565 4201933.129685088  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "104_1"
626131.6740619033 4202440.10714417  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "105_0"
625960.146360933 4202612.8754013805  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "105_1"
625635.5335016225 4202861.385089041  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "105_2"
625467.247181127 4203003.611074079  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "106_0"
625453.2195 4203113.971190821  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "106_1"
625472.3165260282 4203437.908019256  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "106_2"
624664.3072897275 4204562.861579526  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "107_0"
625037.5740154854 4203985.569619767  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "108_0"
625022.7718083062 4204369.119935634  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "108_1"
625497.094352612 4204490.262985547  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "108_2"
624954.989653164 4204855.093088226  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "108_3"
624731.0591006691 4205043.721977405  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "111_0"
624756.4546025555 4205269.783976333  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "111_1"
625176.7272708209 4205616.319444608  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "111_2"
625467.6404835056 4206304.316940054  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "111_3"
625620.7793605478 4206635.506591036  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "114_0"
625486.5412147322 4206483.202199462  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "114_1"
625194.4807819157 4206772.932058473  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "114_2"
624830.7580076044 4206869.759658945  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "115_0"
625533.9483502156 4207295.40415072  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "116_0"
625019.4040735752 4207307.244020643  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "116_1"
624754.128136755 4208333.866949596  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "117_0"
624724.3783121371 4208981.071688506  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "117_1"
624792.8333766848 4209795.027765584  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "117_2"
626322.1293403406 4208711.619207495  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "118_0"
625472.934758171 4208759.484241921  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "118_1"
625745.0924084372 4207872.426781475  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "118_2"
624936.431099843 4207864.485959391  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "118_3"
626381.2452804877 4209450.780593794  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "119_0"
626202.7226498944 4209894.0120070595  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "119_1"
625646.7118257385 4210930.114542504  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "119_2"
625444.3614719992 4211512.011086047  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "119_3"
624799.5132184654 4211417.89662988  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "120_0"
624748.3402797265 4211192.6441845745  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "120_1"
624899.4212814783 4210799.6490042275  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "120_2"
624742.7592071411 4210275.558559777  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "120_3"
624487.5621670119 4210529.382890573  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "121_0"
624375.5990901385 4210985.176689833  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "121_1"
624515.5246052213 4211632.655604595  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "121_2"
624635.4210400245 4212292.069413819  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "122_0"
624587.5149298052 4213019.64488922  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "122_1"
624764.2324846927 4211780.00658487  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "123_0"
624646.1147103403 4212104.43645646  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "123_1"
624824.6766091747 4213614.860124534  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "124_0"
624925.5072611913 4214233.1255290955  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "124_1"
625264.7232544284 4214557.549638019  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "124_2"
642751.8394112618 4187448.1773171537  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "125_0"
642272.8201918973 4188092.525215729  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "125_1"
642153.6145638026 4188575.477075516  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "126_0"
642646.2574515156 4189232.481579141  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "126_1"
642646.3294523031 4189999.0346239163  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "126_2"
642923.854446728 4190869.5139439935  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "127_0"
642952.6388859343 4191426.9405323225  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "127_1"
642699.7074682919 4192627.3356027715  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "128_0"
642825.555374621 4193281.0023116358  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "128_1"
642270.9843852592 4193639.769466811  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "129_0"
641832.2357598671 4194232.682836356  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "129_1"
641300.7195811019 4194474.339000001  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "129_2"
640764.2583590372 4194379.419336226  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "130_0"
639739.7011498791 4194521.865264729  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "130_1"
639425.9697740453 4194704.8116239365  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "130_2"
639021.9185642474 4194899.803368234  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "131_0"
638494.3504008657 4194967.182671037  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "131_1"
637876.5315533702 4194911.077346698  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "131_2"
637346.6316638043 4194753.372591771  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "132_0"
637148.0772269559 4194766.509113861  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "132_1"
636451.8158545722 4194039.0638660146  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "133_0"
636131.4480703415 4193735.116905823  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "133_1"
635389.4883381114 4193981.2212971733  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "133_2"
634364.1003005245 4194287.403600495  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "134_0"
633504.0204189875 4193908.9124021535  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "134_1"
633019.1196389695 4194712.409182516  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "135_0"
632704.1955097571 4195397.858424987  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "135_1"
632354.0176777834 4196058.386469281  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "136_0"
631609.0328317442 4196800.740659211  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "137_0"
631344.3949266709 4196710.532386486  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "137_1"
630950.7012468238 4197173.449106786  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "138_0"
630533.0394600524 4197139.560185384  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "138_1"
630766.4550000001 4197508.699207782  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "139_0"
630601.0767328342 4198100.453328903  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "139_1"
629984.4720377646 4198248.12875907  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "140_0"
629750.1754131834 4198367.8860764755  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "140_1"
629607.4065502759 4198423.392321837  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "140_2"
629535.5955232707 4199168.251538707  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "140_3"
630024.5594691391 4197898.958813331  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "141_0"
629742.1799084187 4198245.385364804  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "141_1"
629473.2320507037 4198512.313795308  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "141_2"
629718.5354818368 4198552.419022981  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "141_3"
629083.7120846291 4198553.236509554  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "142_0"
628974.975766932 4199024.795859034  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "142_1"
629156.0371450894 4199134.1479567615  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "142_2"
629400.1302039617 4199859.306521515  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "143_0"
629047.2296237429 4200340.935369871  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "144_0"
629048.7779381175 4200505.683985721  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "144_1"
628953.5063034808 4200852.069803794  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "144_2"
629512.8722339044 4200790.125725655  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "145_0"
629031.8155921397 4201090.562784124  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "146_0"
629603.3177575304 4201295.001803369  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "146_1"
629595.9220654863 4201776.06813854  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "147_0"
629138.4380508864 4201503.530384621  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "148_0"
629342.8051764063 4202127.326463354  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "148_1"
629077.3402868904 4202514.175966829  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "149_0"
629022.8972932228 4202768.01993207  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "149_1"
628950.3251499485 4203257.900602816  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "149_2"
628548.3002854174 4203807.267715749  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "150_0"
628774.8990169521 4204680.563699202  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "150_1"
629501.4969 4205072.040183536  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "151_0"
629121.3694073143 4205490.268386061  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "152_0"
629254.4375960171 4206135.967776921  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "152_1"
629430.8500886712 4206415.396853038  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "153_0"
629767.0228865733 4206630.047777835  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "153_1"
630214.824141301 4206994.070096641  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "154_0"
630340.0944818355 4206939.482005582  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "154_1"
630785.6289732513 4206696.295155013  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "154_2"
630902.8614747247 4207515.277630321  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "155_0"
630488.1108939154 4207536.932921141  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "156_0"
630314.2614375227 4207994.705760092  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "156_1"
630617.463399898 4208163.170027875  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "157_0"
630673.6591519141 4207644.042173684  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "158_0"
630427.4067722695 4208322.321042298  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "159_0"
630387.1819319759 4208561.831726414  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "159_1"
630500.456904574 4208860.691112189  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "159_2"
630646.6078474444 4209342.861793431  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "160_0"
631345.0758246158 4209582.317096717  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "160_1"
632127.621039214 4209938.837018178  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "160_2"
629788.5425655025 4209557.443200001  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "161_0"
629799.0897110413 4209794.07612263  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "161_1"
630011.2612333933 4210887.872926427  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "161_2"
629676.6938535738 4211722.553877246  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "162_0"
629928.1579884749 4212236.286406846  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "162_1"
630052.2624869662 4212485.838099273  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "162_2"
628752.1492836986 4212079.278841166  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "163_0"
628769.6226171681 4212615.014381446  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "163_1"
630855.433853368 4204192.836322423  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "164_0"
630755.8880249596 4204539.824408518  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "164_1"
630565.8203847047 4204844.010684868  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "165_0"
630375.8157 4205167.103982579  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "165_1"
630466.9749513316 4205298.197579116  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "165_2"
630943.7950878902 4205798.149278989  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "166_0"
631247.9475637208 4206404.541135212  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "167_0"
630885.2642232472 4206974.01792866  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "167_1"
630713.5470999768 4206100.33819758  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "168_0"
630630.7076186985 4206677.599710095  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "168_1"
635728.5853413058 4205975.137869837  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "172_0"
636491.91697556 4206369.044375915  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "172_1"
634356.2160245829 4205085.551882791  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "173_0"
634528.680977969 4205126.018460055  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "173_1"
634971.1353479946 4205419.403121993  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "173_2"
635375.3589833329 4205677.510945204  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "173_3"
634187.2089665256 4203895.552024426  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "174_0"
634169.5069663774 4204018.416104708  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "174_1"
634033.6531785288 4204635.198867566  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "174_2"
634078.3374308003 4204916.281456225  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "174_3"
632656.5579 4203646.152  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "175_0"
632979.6459 4203608.3568  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "175_1"
633549.8505000001 4203627.2544  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "175_2"
631586.2395620771 4203641.8115851935  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "176_0"
632105.416267444 4203627.266459989  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "176_1"
629828.7271406627 4203568.832819127  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "177_0"
630471.4145942922 4203550.515148438  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "177_1"
629168.1727240062 4203003.079381404  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "178_0"
629247.6460664399 4203265.165540997  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "178_1"
629095.596737436 4203402.915040045  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "179_0"
637527.8076964758 4200217.869368979  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "180_0"
636917.742304662 4201169.363894845  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "180_1"
636571.786552879 4201460.035774533  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "180_2"
636144.6954855078 4201702.239641856  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "180_3"
635831.6282141565 4202108.187560362  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "181_0"
635622.3663759567 4202359.218504903  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "181_1"
634888.546622982 4203258.5731720645  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "181_2"
634262.695676026 4202971.261141685  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "182_0"
634060.9546571614 4203192.551601313  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "182_1"
633909.3419708783 4203406.021763321  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "182_2"
639069.7109785796 4184250.26453024  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "183_0"
639259.3823378634 4182917.1252071424  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "184_0"
642916.8805834092 4185596.3011420057  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "199_0"
641884.1059666073 4185823.8389357673  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "199_1"
644689.9185660603 4183596.349274222  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "201_0"
643916.4603675233 4184713.5016257814  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "201_1"
643254.5569490709 4185146.504961798  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "202_0"
641808.9982665995 4185550.0879536183  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "202_1"
641354.9113529318 4185159.5832202905  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "203_0"
639985.3750527801 4185214.863592039  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "203_1"
640112.365025598 4186911.8895244207  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "204_0"
639679.5155592891 4186906.3991186484  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "204_1"
639261.3993861914 4186916.911572716  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "204_2"
638742.6241032258 4186900.884580087  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "204_3"
638360.8446164505 4186810.934379119  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "204_4"
639097.4405628588 4186245.28772188  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "205_0"
638872.8849076281 4186509.3823559107  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "205_1"
638428.048412823 4186931.137054674  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "205_2"
638096.1078293507 4186818.643195862  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "206_0"
637274.2564040847 4186802.1855871947  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "206_1"
636720.8878639108 4186785.7375250184  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "206_2"
636249.7183001669 4186785.7279587314  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "207_0"
635822.3417781462 4186769.2827454293  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "207_1"
635290.8937416598 4186780.2327089924  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "208_0"
634934.7741263221 4186769.244141078  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "208_1"
634474.5244250025 4186736.3482605116  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "208_2"
633953.9663372874 4186714.52454007  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "209_0"
633389.6559930332 4186709.19094878  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "209_1"
632803.4410274414 4187016.0354000004  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "210_0"
632392.5096451172 4187005.0778362793  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "210_1"
631872.0255735954 4186720.1848374745  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "211_0"
631422.7537027602 4186703.72669726  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "211_1"
630935.1486804953 4186703.7143028392  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "211_2"
630266.6894047557 4186665.33618199  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "212_0"
629635.7033295799 4186650.127321237  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "212_1"
629071.4363838859 4186664.092134162  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "212_2"
627806.6958823053 4186594.0363734355  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "213_0"
614925.9908144531 4209184.91769668  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "215_0"
614197.9460507124 4209487.297091753  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "215_1"
613484.180657097 4209023.4336  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "215_2"
628095.8874432065 4188094.6489087245  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "217_0"
629000.7327620257 4189960.9369492433  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "219_0"
628561.9472868455 4189902.551321384  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "221_0"
627731.052743552 4190888.946217211  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "225_0"
632802.6505589202 4194388.7462894125  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "226_0"
630511.500685548 4193126.396185222  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "228_0"
629569.3062863536 4192566.343585162  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "229_0"
628852.5009706717 4192118.5641810223  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "230_0"
626772.2337216382 4190964.7191315684  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "231_0"
627446.8692876499 4188187.2540549147  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "232_0"
630119.9759394232 4197157.472159869  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "233_0"
629480.141948777 4197145.376180806  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "233_1"
628028.0556000001 4197416.04  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "234_0"
627125.9317727293 4196991.942678914  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "235_0"
626604.828867063 4197012.533792926  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "235_1"
625698.2417681586 4197282.142350075  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "236_0"
624936.9096518847 4197533.117897694  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "237_0"
624437.5613305786 4197839.082219396  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "237_1"
623961.3465622131 4197665.97100343  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "238_0"
623495.5764495697 4197488.646957665  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "238_1"
622874.787879914 4197399.611749572  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "238_2"
622574.761581245 4198164.225707107  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "239_0"
622472.5168857588 4199344.356965786  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "240_0"
622549.8350186907 4200295.094435205  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "241_0"
622456.1907892897 4201044.4672023915  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "241_1"
622810.0939314937 4202207.414951003  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "242_0"
623557.1699444035 4203178.52773539  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "243_0"
624030.6549423418 4203345.140975534  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "244_0"
623056.6152 4203967.4112  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "245_0"
621939.0492859777 4203994.354812962  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "246_0"
620322.5160731828 4204091.181195081  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "247_0"
629294.4672419676 4207444.507777393  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "248_0"
628947.8704971046 4207474.344173665  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "248_1"
628352.0421380441 4207772.453332703  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "249_0"
627849.1181668479 4208159.539747124  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "249_1"
627284.6804342131 4208170.564275341  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "249_2"
626631.75730301 4207694.584784966  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "250_0"
626555.4543239629 4207466.405431943  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "250_1"
626099.6155827983 4207105.5535279345  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "250_2"
627045.8302846176 4208194.652034572  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "251_0"
626863.834930469 4208507.56173081  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "251_1"
623495.761126118 4188718.330520668  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "252_0"
624084.3536518387 4189796.6824608627  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "253_0"
624664.8901865748 4190821.7203198327  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "254_0"
625066.3761817936 4191210.5310581033  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "255_0"
625622.8714454776 4190760.9534169864  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "255_1"
625286.2553406077 4191514.2715017386  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "257_0"
628710.8720397841 4200042.875823079  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "258_0"
626715.2439 4200361.6272  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "259_0"
612931.2799996024 4209133.906192228  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "260_0"
612358.0674867758 4209285.845843007  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "260_1"
612120.7376790438 4209407.429288802  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "260_2"
621125.3030943967 4204584.625079141  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "261_0"
621056.2204186663 4205872.866313246  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "261_1"
621241.4857999057 4207267.736625929  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "262_0"
621365.1219959927 4207725.444310347  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "262_1"
620764.9165902773 4206712.232549797  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "263_0"
620601.3228495115 4207219.4111826345  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "263_1"
622783.7382230833 4208843.642288078  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "264_0"
623592.0358616703 4209537.626181848  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "264_1"
622329.5477499817 4208488.1869303575  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "265_0"
621930.3059741168 4208206.567616567  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "265_1"
620996.8057161327 4207501.776844425  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "266_0"
620714.9377711598 4207559.901103895  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "266_1"
620899.5411638547 4207875.645262453  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "267_0"
622101.383404618 4209494.095069745  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "268_0"
621803.0985175847 4209931.792030099  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "268_1"
621534.9533762411 4210229.034587547  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "268_2"
621340.0814984374 4210490.140469557  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "268_3"
620497.4203966673 4211002.424919873  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "269_0"
619969.844693604 4211537.948725317  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "269_1"
619394.2901477696 4211943.881603493  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "269_2"
618391.8128386582 4211937.451132704  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "269_3"
618248.8421142655 4212029.6531939935  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "270_0"
617981.8433419478 4212267.322682192  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "270_1"
617812.5397611579 4212418.265209602  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "270_2"
617849.706005697 4212565.488735343  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "270_3"
617948.4177188481 4212704.915963206  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "270_4"
618617.9037838562 4208707.960250878  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "271_0"
617860.2514825976 4209203.472448895  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "271_1"
616837.4425184027 4210141.175049896  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "271_2"
616630.6375814105 4210593.213218725  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "272_0"
616823.6249981702 4211165.5973398695  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "272_1"
617936.1798666518 4211950.107928249  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "272_2"
619751.918301256 4208078.170635617  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "273_0"
618534.3666093267 4207934.637727015  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "274_0"
616793.6074667438 4207938.245023514  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "274_1"
615835.5960778499 4208113.841840245  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "274_2"
615178.2472069854 4208906.6857677465  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "275_0"
614772.5303280927 4209674.121151062  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "275_1"
612867.0311906396 4209317.95160589  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "275_2"
612126.5040498379 4209531.209545248  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "275_3"
623988.8778795874 4213984.848826258  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "276_0"
623398.4948277173 4214036.205837684  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "276_1"
622892.0608977469 4213620.861101485  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "276_2"
622722.6680098159 4213119.1655199  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "276_3"
621974.493527677 4213775.926557141  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "277_0"
621689.6610618959 4213949.0601232  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "277_1"
620929.8200960272 4213035.780781898  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "277_2"
620625.6998220644 4212408.4711741125  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "277_3"
620031.2886636681 4212419.889960543  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "278_0"
619937.7459453827 4212538.083060704  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "278_1"
619586.2133168471 4212856.173946085  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "278_2"
619178.6957843335 4212972.313627508  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "278_3"
618849.8144400849 4213020.460447552  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "278_4"
618503.5748517233 4212687.126487917  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "279_0"
618177.1230938948 4212949.831404166  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "279_1"
617845.090093532 4213196.181042479  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "279_2"
617186.9816582204 4213101.749054883  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "279_3"
616614.9067637797 4213250.655798294  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "279_4"
607027.2907137921 4210785.644208618  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "283_0"
607728.5498005819 4210304.594153928  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "283_1"
608020.704892627 4209967.914180567  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "283_2"
608306.2991954543 4209893.1919749025  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "284_0"
607937.9615954087 4209478.712948197  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "284_1"
607465.836980795 4209345.810618799  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "284_2"
607007.4509866635 4209196.461817082  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "284_3"
602400.418716965 4211786.577891008  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "285_0"
602501.6611402073 4211513.6116503775  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "285_1"
602517.4824352985 4211159.998890675  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "285_2"
602619.5016290057 4210848.013079981  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "285_3"
602815.9043334333 4210339.42633688  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "285_4"
603038.1414958263 4210134.147773298  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "285_5"
602285.3737022602 4212958.139534248  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "286_0"
602364.8623700589 4212715.590217248  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "286_1"
602502.174286277 4212323.519735284  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "286_2"
602455.6604447208 4212112.1310424395  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "286_3"
602478.2005329079 4209314.447205806  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "287_0"
602231.2366037547 4209190.563899681  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "287_1"
601877.4484674025 4209178.018703742  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "287_2"
601509.8746686765 4209693.432384551  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "287_3"
601159.9710303701 4209883.082136057  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "287_4"
600346.56850932 4209679.950711345  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "288_0"
599940.9390951529 4210084.639314219  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "288_1"
599580.5908679798 4210170.872071174  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "288_2"
599277.0342187006 4210250.497593661  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "288_3"
598945.3883366673 4210376.673157713  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "288_4"
598689.722047023 4210566.568971823  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "288_5"
598481.8007198247 4210730.900212727  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "288_6"
601082.7773262803 4210823.738958249  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "289_0"
600767.475773118 4211282.07053696  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "289_1"
600447.8670018978 4211598.827209691  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "289_2"
600386.1376259741 4213146.725698586  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "290_0"
599792.1914725193 4212632.155435878  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "290_1"
599245.3578036304 4212205.375591096  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "290_2"
598919.7322441615 4211926.373675132  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "291_0"
598171.894051239 4211472.652037089  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "291_1"
600269.9115505092 4212186.254162917  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "292_0"
600269.8756662521 4212382.661889337  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "292_1"
600597.1089322998 4212791.625710941  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "292_2"
599532.8089449572 4212102.144560572  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "293_0"
599759.8086221908 4211982.118350495  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "293_1"
599970.1237376117 4211914.612000395  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "293_2"
600108.4509617665 4211888.141233672  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "293_3"
599567.5260761724 4211840.998612382  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "294_0"
599375.5779555517 4211504.502864969  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "294_1"
599135.5000121847 4211329.543991434  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "294_2"
598568.3322736968 4211046.0341763655  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "294_3"
606755.8396644692 4210677.88025232  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "299_0"
606776.2173524213 4210341.539549441  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "299_1"
606776.225924774 4209883.898642655  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "299_2"
606746.0305009496 4209550.564084852  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "299_3"
606526.6144835263 4209139.684163942  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "300_0"
605931.0864375802 4208956.385356285  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "300_1"
605198.095617999 4208841.65132308  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "300_2"
615097.0564993464 4219147.277135597  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "309_0"
614901.7311707779 4218954.393379884  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "309_1"
614771.054288644 4218745.434664651  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "309_2"
614666.8049798699 4218406.260666555  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "309_3"
614405.7962692293 4218171.255670554  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "309_4"
614166.478391441 4218561.080051526  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "309_5"
615509.7992404248 4216665.217502544  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "310_0"
615397.5642179878 4216891.947747842  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "310_1"
615397.5174209581 4217180.07943887  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "310_2"
615454.3773750998 4217459.826011046  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "310_3"
615592.5121542416 4217729.317435835  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "310_4"
615423.6836730907 4218067.696681428  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "310_5"
615501.8656863996 4218353.7461612  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "310_6"
615554.0835862746 4218667.225570594  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "310_7"
615645.4352212271 4219001.265774017  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "310_8"
641812.3129283366 4208821.4276065435  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "311_0"
640843.5644236852 4209937.2375426935  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "311_1"
640108.3693718553 4211144.484617539  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "311_2"
639408.0130870498 4212010.787698857  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "311_3"
641714.3863214045 4208049.006285126  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "312_0"
640972.7971754938 4207554.579135519  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "312_1"
639247.2762256952 4206607.95435887  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "312_2"
638110.2204828808 4211458.1049337  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "313_0"
637450.5577651245 4211329.40722078  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "313_1"
636586.3799693282 4211995.130993952  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "313_2"
635573.098857166 4212960.665538492  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "313_3"
634711.6973749335 4212315.195209503  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "314_0"
633490.9864959317 4211367.0182102425  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "314_1"
633646.5012892266 4211215.7987114675  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "315_0"
634338.5148117673 4210260.559584204  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "315_1"
632970.565450883 4210989.666020402  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "316_0"
639168.4527801911 4215870.284479715  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "317_0"
639068.6559226239 4214930.551713084  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "317_1"
639168.1861255363 4212174.498157455  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "317_2"
635320.5206776023 4213814.045201962  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "318_0"
631731.6595467287 4214141.794834565  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "319_0"
631819.8612468536 4213233.061878388  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "319_1"
638161.4405856688 4216121.148918498  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "320_0"
637136.4215440801 4215799.345499995  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "320_1"
636654.1743554802 4215632.721856645  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "320_2"
635344.4111380501 4214482.690847974  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "320_3"
634323.7270131565 4216176.863395008  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "321_0"
634490.9857931557 4215934.463961794  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "321_1"
634988.1141501458 4214990.682675114  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "321_2"
635210.5091954725 4214589.278826394  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "321_3"
632515.6970763712 4217140.024435799  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "322_0"
633300.7473019382 4217004.005648891  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "322_1"
633890.7755327981 4216741.752791847  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "322_2"
631829.9098274414 4219401.095285045  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "323_0"
631762.3836360396 4218959.782397053  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "323_1"
632036.8809569423 4218780.917446057  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "323_2"
632543.2485 4218416.455220796  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "324_0"
632360.5894489576 4217941.546265546  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "324_1"
632324.0060953286 4217466.287430587  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "324_2"
632031.6012198412 4217478.513977935  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "325_0"
631593.4002723648 4217064.659585456  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "325_1"
631276.6572196713 4215968.607863221  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "325_2"
631216.3994213176 4215072.09201484  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "326_0"
630194.772021737 4216613.02816848  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "326_1"
629473.8057865291 4216971.338439952  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "327_0"
628810.6626829918 4216696.42599927  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "327_1"
627951.8879856372 4216488.307351131  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "327_2"
627046.6871268951 4216176.673186894  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "328_0"
626490.8062954514 4215826.49592861  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "328_1"
625893.7726144762 4216114.582596982  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "328_2"
631593.3902522699 4235369.095203491  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "329_0"
631807.4819199716 4234427.841258227  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "330_0"
632011.3653707419 4233686.232844788  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "331_0"
631778.422124079 4233271.246213455  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "331_1"
631699.8466292804 4233157.741783136  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "331_2"
631138.0587971812 4232627.823012132  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "332_0"
630668.0011897056 4232337.180586895  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "332_1"
630734.80273821 4232071.654713101  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "332_2"
631759.4785099928 4232768.024845681  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "333_0"
635689.6041648106 4235371.102917392  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "334_0"
634007.8213440272 4236002.566523741  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "334_1"
632767.9127948716 4233593.50916321  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "335_0"
632167.5206854431 4232417.796631495  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "336_0"
631831.7640991658 4231396.843098698  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "337_0"
631590.959786683 4230870.075834317  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "337_1"
631801.5984450905 4230620.347922539  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "337_2"
633338.1334054 4229521.514530012  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "338_0"
633440.0606935369 4229380.784651089  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "338_1"
632919.4831713332 4227894.027750716  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "339_0"
632565.3909129568 4227333.63003965  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "339_1"
631767.3832908992 4226489.604379859  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "340_0"
631794.775117636 4226059.219933362  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "340_1"
631916.9328962932 4224839.317571839  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "341_0"
631760.2381089454 4224806.321223799  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "341_1"
631297.485030442 4223916.340614378  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "341_2"
631017.0377211071 4223090.7167652575  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "342_0"
631199.531327769 4222739.149197731  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "342_1"
631060.2827829922 4221690.320125105  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "343_0"
631356.9734840404 4221519.915507551  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "343_1"
631597.0834543802 4221391.681988149  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "344_0"
632177.8930506728 4219804.8017460415  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "344_1"
631569.0170723766 4219573.430386845  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "345_0"
630967.2924211777 4220105.455911002  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "345_1"
629810.5822145301 4220126.887401454  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "345_2"
628559.9962611014 4219840.716654068  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "346_0"
627245.4040565013 4219600.3858342655  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "346_1"
626447.8337376429 4220195.683768922  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "347_0"
626127.1024558957 4221326.743080848  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "347_1"
624298.2146286584 4219901.864234116  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "348_0"
624307.4915362793 4219570.962481945  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "348_1"
624753.0526371283 4219341.068336528  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "349_0"
625540.5074641806 4219045.1624792935  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "349_1"
626332.1484000001 4217936.055812904  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "349_2"
625937.3084500184 4217077.6842597835  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "349_3"
635848.396774292 4229423.353403121  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "350_0"
634302.0823990433 4228163.684805908  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "351_0"
633349.5188662752 4228713.468621063  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "351_1"
635851.1739253559 4225547.605543443  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "352_0"
634851.795777869 4225403.551423938  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "352_1"
634031.6296754607 4225296.634020095  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "353_0"
633290.0218889263 4224887.554393926  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "353_1"
632343.2264081378 4225775.779859122  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "353_2"
636537.4508127914 4222578.163324703  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "354_0"
635772.9668106475 4221691.320863168  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "354_1"
635179.3027264001 4222871.862311057  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "354_2"
631797.5304173324 4222440.527145968  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "355_0"
631317.8193365326 4222153.703949306  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "355_1"
631433.5700619061 4232086.639201681  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "356_0"
630822.9945570943 4231701.064876077  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "356_1"
630849.1885511195 4231148.191715064  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "357_0"
630595.6939082539 4229540.272172047  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "358_0"
630408.3281654352 4229337.621088948  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "358_1"
629775.7929369193 4229477.130692674  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "359_0"
629266.6616329813 4228741.17209239  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "360_0"
628951.7959541873 4228569.3858670965  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "360_1"
629234.4309087924 4227582.246131766  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "360_2"
629252.587955382 4226607.502250877  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "361_0"
628929.4804360616 4225342.316833806  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "362_0"
628510.4675869404 4223930.907858107  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "362_1"
628417.7113225596 4223674.873312553  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "362_2"
627819.2613173987 4223306.665211773  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "362_3"
627795.2163997155 4223263.621399894  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "362_4"
627149.7319863514 4222949.044562151  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "363_0"
626620.7710568954 4222735.8383658845  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "363_1"
626463.2052333748 4222448.302258042  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "364_0"
625881.7434570069 4221664.992671364  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "364_1"
630796.3842841868 4234302.380657206  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "365_0"
630999.1736201756 4234249.920397619  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "365_1"
631199.3064772546 4234201.161287963  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "365_2"
629851.3785559447 4233201.291164494  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "366_0"
629445.2857779714 4232494.498275073  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "366_1"
627625.867997973 4230960.686666427  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "368_0"
627772.689298416 4231038.721326283  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "368_1"
627843.4880473664 4229605.969451632  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "369_0"
626939.3742981296 4228216.670995968  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "369_1"
626317.0283317596 4227602.34170347  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "370_0"
625185.4532411563 4226850.302710145  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "370_1"
624615.4994894487 4226059.69144065  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "371_0"
624062.2425479245 4224306.493934832  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "372_0"
623584.8910294754 4223724.358252264  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "372_1"
622815.0603882615 4222994.845554253  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "373_0"
623419.9188092089 4221804.018808104  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "374_0"
623945.1735848145 4220980.006072558  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "374_1"
624481.0119941195 4221062.119200001  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "374_2"
624944.8096807491 4246060.831186895  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "377_0"
624064.3474420664 4243726.9640220795  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "378_0"
624513.4431023239 4243285.836044594  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "379_0"
624234.1913306725 4243422.82180233  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "379_1"
624025.4676982482 4243657.7697076555  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "379_2"
623910.228138441 4243505.423129615  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "380_0"
623698.9333682489 4243213.827459266  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "380_1"
623384.8120921886 4242528.4716761885  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "380_2"
623482.6488292324 4242157.533816332  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "380_3"
623102.0837315496 4241517.721474582  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "380_4"
622540.5536113421 4240404.153049879  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "381_0"
622069.8774868045 4239565.222967644  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "381_1"
622386.393602311 4238803.840729573  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "381_2"
622110.3012125007 4238506.245133331  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "381_3"
622079.158487941 4238444.854491141  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "382_0"
622532.5751806549 4237999.811723651  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "382_1"
622605.615252543 4237415.192769498  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "382_2"
622220.7165198823 4236934.314475718  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "382_3"
622321.0735314309 4236397.350072434  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "382_4"
622515.8200410914 4235040.1540012555  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "382_5"
624693.2369071438 4240485.973200616  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "383_0"
624263.6760887206 4240124.697637205  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "383_1"
624213.1814391501 4238840.411290181  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "383_2"
623560.6450809037 4238191.392446768  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "383_3"
623609.0462774163 4237857.245440112  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "383_4"
623620.7385295782 4236404.776572016  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "384_0"
623147.2338213098 4235655.479702815  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "384_1"
622564.802751414 4235117.35638997  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "384_2"
622525.6911904238 4233515.857192607  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "385_0"
622537.5586255628 4232684.431123687  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "385_1"
622549.4390149325 4231556.029372574  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "386_0"
622190.3788700665 4230350.011605108  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "386_1"
621836.7367643485 4229905.0630554315  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "386_2"
621911.3790163412 4229486.959532089  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "386_3"
621692.1480489657 4228682.974705057  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "386_4"
620969.7369983646 4228111.666659118  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "386_5"
620023.9016641901 4228009.482979521  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "387_0"
619463.5059088337 4227879.237039241  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "387_1"
619061.5985905783 4227586.976876356  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "387_2"
618842.455978274 4227294.722182065  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "387_3"
618526.0482943455 4227098.096680261  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "387_4"
617590.8504893894 4226660.190400908  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "387_5"
621838.3296 4238671.3296  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "388_0"
621341.6291344517 4238633.836462717  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "388_1"
621180.7584997425 4239132.563914671  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "388_2"
620397.1351737734 4238866.366125217  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "388_3"
619366.6074056679 4238878.428737064  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "388_4"
618563.2041778011 4238662.529752713  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "389_0"
619170.3522423415 4237634.27301167  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "389_1"
618659.7687801453 4235953.67003016  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "390_0"
618042.9600000001 4235113.399272232  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "390_1"
617862.4663908087 4234836.751399073  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "390_2"
617450.186608575 4234023.603505422  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "390_3"
617061.5849504527 4233408.571950871  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "390_4"
623799.4926157537 4267642.4139284035  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "391_0"
623536.9519099568 4266958.787362887  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "391_1"
623660.6518181919 4265258.165174171  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "392_0"
623724.7317466412 4260562.768885819  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "392_1"
623682.0022902444 4258575.223014481  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "393_0"
622420.9964499259 4255005.746799603  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "393_1"
621772.0932264293 4253326.107602055  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "394_0"
620829.6615233434 4250085.507671849  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "394_1"
619656.8329510391 4247402.236518479  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "395_0"
618885.0848861212 4244940.068798351  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "395_1"
618297.1683277205 4243029.228856883  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "396_0"
618071.044098496 4241150.375837002  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "396_1"
617709.1907113924 4239115.438715438  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "396_2"
616339.8519 4231971.216  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "398_0"
616498.8565106023 4231272.759620198  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "398_1"
617264.3374467677 4230200.236724747  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "398_2"
617782.9200205804 4229815.58397447  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "398_3"
617819.3892 4228719.595351322  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "398_4"
617999.0726653113 4228047.353322344  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "398_5"
617673.2387613528 4227513.82384666  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "398_6"
617490.5126723201 4227038.949504358  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "398_7"
616791.4294173252 4243649.3234346695  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "399_0"
616954.0623968729 4241349.721635487  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "399_1"
616876.7710240964 4238913.246946298  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "399_2"
616905.9757028578 4237363.543702555  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "400_0"
616467.5272155008 4236048.445306594  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "400_1"
615766.0201163037 4233651.796007555  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "400_2"
614480.0072123867 4241530.826809621  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "401_0"
614610.3362459465 4238872.092174785  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "401_1"
614427.6278298349 4237165.586036533  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "401_2"
612025.1948587243 4238596.264482324  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "402_0"
613281.5857962095 4237364.055481566  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "402_1"
614012.3602692469 4236341.116049462  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "402_2"
614830.7871377375 4235171.7684110245  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "403_0"
615093.8548192304 4234060.395315162  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "403_1"
614973.6582126687 4233768.011570956  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "404_0"
615241.6601022616 4233481.736458848  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "404_1"
615290.175044287 4233276.645599301  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "404_2"
615672.9471400644 4232926.035895274  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "405_0"
611264.8661943448 4234996.600357537  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "408_0"
611690.8046876638 4234956.862337226  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "408_1"
611944.7483880486 4234515.11703855  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "409_0"
613219.9837793793 4234402.429960087  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "409_1"
614450.8700786096 4233535.040986712  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "409_2"
630289.6556956437 4271766.474296901  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "410_0"
629986.1222241328 4270553.111842863  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "410_1"
629162.3685358001 4269675.640952499  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "410_2"
629609.2175020601 4268709.80230912  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "411_0"
629931.1583348142 4266999.054325714  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "411_1"
628445.7412408069 4265455.896973533  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "411_2"
627597.8745190622 4264046.733184211  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "412_0"
626366.9138621266 4263618.978324976  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "412_1"
626068.9763501649 4262599.957812672  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "412_2"
626065.2178276688 4261982.818304263  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "413_0"
626290.9184491688 4261651.313474038  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "413_1"
627027.8366797192 4260145.829074516  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "413_2"
627875.2191154322 4259790.799522758  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "413_3"
628816.733560955 4259154.024777641  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "414_0"
630305.7025704266 4259504.10801292  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "414_1"
630826.3082743565 4258934.562531536  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "414_2"
630897.7049125001 4257494.247342492  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "414_3"
631018.9373947647 4256393.799734822  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "414_4"
630375.3499651671 4255283.996178517  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "415_0"
629255.1532385362 4254879.451775142  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "415_1"
628504.510874509 4255313.363872559  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "415_2"
628398.4760953177 4254332.682635318  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "415_3"
629182.2516993716 4253239.403997375  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "416_0"
629693.6703923226 4252358.391694883  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "416_1"
630066.6575147071 4250885.770154044  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "416_2"
630066.6668605797 4250166.2408018075  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "416_3"
629162.3650066456 4248330.169382832  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "417_0"
629469.1483194598 4247550.600205475  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "417_1"
626002.3846797416 4244759.645661649  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "418_0"
625273.4201816454 4243889.554502303  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "418_1"
624749.6656505851 4243041.044489769  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "418_2"
624697.7705735305 4242923.032560428  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "419_0"
624476.1187137775 4241972.999514975  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "419_1"
624930.0152054367 4240864.536493637  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "419_2"
625034.9900993651 4240603.280314626  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "420_0"
626362.8377704691 4238835.990411478  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "420_1"
628343.7531238582 4237035.5512930155  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "421_0"
629547.4752864469 4235953.747179083  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "421_1"
630385.0563991799 4235035.352865309  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "421_2"
630483.0624995133 4234363.129535981  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "421_3"
630247.3106822227 4233837.242821652  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "422_0"
629953.6958417243 4233391.254419406  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "422_1"
629583.7624729079 4233282.646953927  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "423_0"
627342.7982101076 4233750.2574000005  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "423_1"
626498.4179016647 4232217.618935729  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "424_0"
626581.08165551 4229575.881938737  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "424_1"
626295.8574172651 4228746.115862278  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "426_0"
625431.4889234065 4228020.058223356  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "426_1"
624352.3204354658 4227209.4753356725  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "427_0"
623774.0400442358 4226292.264411272  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "427_1"
622381.5316494522 4224810.023529311  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "427_2"
621359.8277836248 4225037.3316738745  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "428_0"
620362.0824753598 4225481.632936872  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "428_1"
618989.5770008505 4225749.522972342  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "429_0"
618091.0094945444 4226226.6789444545  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "429_1"
617606.2753613348 4226297.5325265  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "429_2"
616956.7860207078 4226556.638522476  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "429_3"
616796.205092581 4225650.510774375  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "430_0"
616538.8918794041 4225368.942020182  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "430_1"
616426.367147709 4224618.890856855  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "430_2"
615956.099563313 4224079.692021295  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "430_3"
615685.6837846689 4223737.563820741  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "430_4"
615404.3953519245 4222903.196918784  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "430_5"
615334.9178297117 4222216.152754208  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "431_0"
615188.6940287314 4221576.768332283  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "431_1"
614932.9805432698 4220498.83050368  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "431_2"
614439.5539699054 4219402.723527779  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "431_3"
613964.6037905473 4218800.201071087  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "431_4"
613615.8888580413 4217108.494133202  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "432_0"
613148.2730135429 4215879.553679327  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "432_1"
611491.5415528445 4215399.978913396  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "432_2"
612886.83538212 4217868.71601346  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "433_0"
612409.9169999429 4216940.199290349  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "433_1"
611278.0223882376 4216335.990354512  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "433_2"
610075.8449529399 4215373.529685899  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "434_0"
608397.130860817 4214187.913470031  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "434_1"
606604.7526543139 4212972.878076204  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "434_2"
605425.4877282652 4212570.724893224  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "435_0"
604710.5973879158 4213696.40276215  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "435_1"
604166.63748582 4214031.79794024  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "435_2"
603155.0288753387 4214246.5005375305  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "435_3"
602563.8867553456 4214553.4494737135  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "436_0"
602125.2027084155 4214697.215443605  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "436_1"
601578.2515734263 4214960.830659778  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "436_2"
601171.591333857 4213335.795000855  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "436_3"
600876.7468711964 4213186.749868104  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "436_4"
597448.7375472697 4210767.813454109  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "437_0"
596296.809438017 4212233.003167746  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "437_1"
595433.6667596261 4212072.989880315  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "437_2"
594282.6041835522 4212296.917221525  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "437_3"
593724.416224454 4212208.698022457  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "437_4"
593017.6005453145 4212652.854057393  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "437_5"
588598.393235147 4213186.037360835  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "438_0"
587458.7186447561 4213595.582572383  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "438_1"
586357.1644096528 4213786.97160936  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "438_2"
585101.5009939661 4212575.844267034  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "438_3"
584401.590269261 4213973.59916724  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "439_0"
583375.8681636045 4212285.72285876  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "439_1"
582199.8758428671 4212041.6067092875  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "439_2"
580901.9530519216 4211064.100817923  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "440_0"
579771.7851383897 4211003.148229081  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "440_1"
578840.4828739483 4210773.85719583  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "440_2"
578142.048334532 4209374.402340103  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "441_0"
577114.8151484139 4209353.8093527015  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "441_1"
576140.3303528765 4209113.57863378  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "441_2"
597032.5934531102 4212731.975017485  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "442_0"
596218.4385491664 4213036.756803107  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "442_1"
595696.5110373334 4213828.315626884  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "442_2"
592248.1987700439 4211842.63754246  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "443_0"
591240.363267514 4211460.960846143  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "443_1"
590469.5950897379 4213068.808271531  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "443_2"
589482.3112464823 4213021.929458098  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "443_3"
590110.3181270729 4213186.3661518  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "444_0"
588795.7059774136 4214017.579013143  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "444_1"
587740.9256311659 4214412.954863229  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "444_2"
587075.5178987648 4214560.932876927  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "444_3"
586261.9868563879 4214675.587436618  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "445_0"
585810.0238729876 4215367.729085378  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "445_1"
584796.0652321278 4214637.448903978  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "445_2"
588080.7757506642 4216083.717864441  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "447_0"
586924.7948905802 4216663.829353358  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "447_1"
585977.9551643606 4217312.997849664  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "447_2"
585493.7131290361 4217866.488311186  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "448_0"
584669.2658493832 4218624.610580331  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "448_1"
583491.6976249431 4218669.322444815  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "448_2"
583238.3788788278 4220364.628788139  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "449_0"
583467.4473590773 4219448.132361522  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "449_1"
583391.1630092622 4218500.606253417  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "449_2"
588766.4067340356 4215461.714472873  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "450_0"
589794.4365989293 4215163.368353823  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "450_1"
590108.3500826264 4214847.907836876  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "450_2"
582688.5650347274 4217035.085616239  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "451_0"
581955.6094885853 4216256.311477993  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "451_1"
580962.9660448893 4215156.622959883  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "451_2"
584536.4256539899 4212499.643869617  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "452_0"
583223.1672698999 4211919.29351399  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "452_1"
581883.3248755786 4212864.074017742  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "452_2"
584505.1482929413 4215952.120383624  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "453_0"
583100.9544070817 4214405.107319974  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "453_1"
582394.8306229493 4214321.129232633  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "453_2"
582077.6091940238 4213372.582780174  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "453_3"
580092.6934498876 4213415.944355231  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "454_0"
579023.6252633064 4212530.1640351545  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "454_1"
578214.4333865975 4211820.020271027  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "454_2"
584818.0292084396 4230216.983123659  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "459_0"
584676.0431719295 4229358.362871551  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "460_0"
584202.1524719589 4228426.214857288  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "460_1"
583673.7490596302 4227283.626173904  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "461_0"
583026.6279821233 4226981.156846887  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "461_1"
583318.2359004734 4226436.81977225  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "461_2"
582703.0669068597 4225834.770162303  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "462_0"
582287.5124361845 4225476.374467994  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "462_1"
581820.5932878092 4224867.008726703  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "463_0"
582468.8161818461 4224317.78598584  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "463_1"
581611.8486200046 4222950.019601527  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "464_0"
581723.4957741929 4222152.669375705  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "464_1"
580925.0066464185 4221420.62531246  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "464_2"
580623.5664306 4220621.7622405505  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "465_0"
580951.7978902244 4219996.161083544  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "465_1"
581984.2606611325 4219994.795475748  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "466_0"
577851.0001503599 4227666.210442609  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "468_0"
578361.5661451172 4227362.130375521  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "468_1"
577666.4564047916 4227013.456227239  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "468_2"
577314.6348465134 4226286.57374098  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "468_3"
577636.4083354373 4225073.809489533  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "468_4"
577720.3245418812 4223620.24452346  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "469_0"
580065.441342826 4223116.883622868  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "470_0"
580163.8785499418 4222685.408846642  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "470_1"
579298.0655459873 4221594.485089731  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "470_2"
579724.0763239212 4220514.404169697  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "471_0"
578946.277336128 4215750.346338618  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "472_0"
579312.4401008413 4216265.67147565  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "472_1"
579713.6456090139 4217828.0337265  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "472_2"
579034.5167033968 4218343.54459185  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "472_3"
578668.0150030615 4215169.864084994  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "473_0"
578542.1594879652 4215261.796881619  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "473_1"
578445.9821562788 4215344.354768761  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "473_2"
578425.3132694977 4215387.382521683  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "473_3"
578940.315370139 4215325.092551246  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "473_4"
578965.4898166249 4223577.778217083  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "474_0"
579879.3120757533 4223155.882018449  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "474_1"
581414.9177589009 4226048.063692048  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "478_0"
582003.6957750553 4225456.433446781  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "478_1"
578756.1567247304 4224730.546801727  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "480_0"
580112.1802363123 4224700.801704584  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "480_1"
579137.7005182263 4224073.4465013025  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "480_2"
578112.2802366876 4224699.336283389  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "481_0"
584272.7529573621 4229359.859524124  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "484_0"
584154.5469911888 4229430.050305298  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "484_1"
583660.9214332685 4229760.522894204  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "484_2"
586124.9005035063 4231442.554030558  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "486_0"
585778.8628776132 4231600.175713003  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "486_1"
585599.089033551 4231386.21718311  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "486_2"
585662.3011744256 4231008.042628976  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "486_3"
584955.063312536 4230721.539752388  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "486_4"
582194.8984499307 4228905.742715347  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "487_0"
583021.7484981505 4229606.27827341  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "487_1"
587356.4228093628 4226942.59770315  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "491_0"
588271.9944709778 4227561.1806244245  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "491_1"
594246.3794458945 4230104.318983918  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "497_0"
594314.5413750984 4229843.010485506  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "497_1"
594273.1777862702 4229631.063284564  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "497_2"
594349.615038947 4229450.399301076  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "497_3"
594514.599695345 4228990.265652653  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "497_4"
594525.9696381572 4228855.451679296  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "497_5"
594406.692664621 4228099.907405434  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "498_0"
594063.6856232375 4227929.059138572  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "498_1"
593821.6774818604 4227525.274792951  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "498_2"
594138.67727751 4226776.036398745  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "498_3"
594610.1698223667 4226473.623463076  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "498_4"
594557.1741770864 4225802.609374943  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "499_0"
594106.815005591 4225666.067465542  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "499_1"
593461.5060570139 4224971.582530711  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "499_2"
579214.5032176758 4219057.580463375  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "500_0"
579006.8602266955 4219926.829345227  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "501_0"
578896.6752295732 4220158.2410553275  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "501_1"
595230.6021489234 4228122.454249666  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "503_0"
595713.8793568638 4227438.447272197  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "503_1"
595869.9651359266 4226440.645371749  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "503_2"
586904.9803796281 4231355.652399438  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "508_0"
586419.9341474461 4231428.482942294  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "508_1"
599619.2861891779 4214187.112563068  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "511_0"
598428.4073810863 4214638.658191875  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "511_1"
598121.1071028035 4214823.431238869  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "511_2"
597984.1011759861 4216402.392025927  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "512_0"
597200.0211550092 4217104.345415934  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "513_0"
597252.0904369315 4217594.701041372  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "513_1"
597352.393615054 4218835.367367205  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "513_2"
597782.835807727 4219790.647633359  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "513_3"
596460.3581979489 4219926.004710752  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "513_4"
595755.4539010476 4220147.177798973  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "513_5"
595249.9615806835 4221056.08395221  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "513_6"
595712.4424970223 4221947.5588963  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "515_0"
595248.9320092808 4222891.343843858  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "515_1"
595278.2060809645 4222971.256523765  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "515_2"
594872.845119743 4223177.308047385  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "515_3"
594892.3257475102 4223264.709497842  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "515_4"
593722.8145197157 4224520.490051644  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "515_5"
593778.3782939406 4224609.760897674  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "515_6"
592952.675802247 4224728.087066606  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "516_0"
592503.9560346558 4225445.857563534  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "516_1"
591748.2207869672 4225490.362215519  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "516_2"
591111.6239945695 4225839.462544677  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "517_0"
590868.6012996704 4226972.210959576  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "517_1"
589713.152895637 4227488.10198234  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "517_2"
588239.1706287583 4226268.469094845  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "522_0"
587337.329043948 4225900.448648726  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "522_1"
586241.1985032033 4225300.121172306  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "522_2"
584916.934528741 4225396.714127391  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "522_3"
584179.619180544 4224470.743459063  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "522_4"
583258.5664117389 4222996.01564124  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "523_0"
582586.7355756321 4221812.632493116  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "523_1"
587390.5241919168 4225061.095215666  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "527_0"
588015.0328613148 4225997.94892537  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "527_1"
582644.4282467632 4223794.039474562  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "528_0"
582865.6739923883 4223689.811911544  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "528_1"
582106.1628901501 4223778.954  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "543_0"
581181.5210818282 4223840.907793387  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "544_0"
581370.5596044029 4223826.031491982  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "544_1"
637023.5291396789 4235408.780169235  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "549_0"
637057.0308761015 4235044.617537773  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "550_0"
635555.368760598 4237665.992724086  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "552_0"
635551.2740166169 4237310.372401309  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "552_1"
633917.1998345192 4236433.597764171  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "553_0"
632391.1888369685 4236143.2516384665  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "553_1"
630538.4042832294 4240868.514772035  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "555_0"
630673.0262097657 4240580.592115994  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "556_0"
631279.794254659 4238948.294264402  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "557_0"
631826.4426902344 4237472.47177407  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "557_1"
631513.8612147486 4236716.49781353  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "558_0"
631494.7174523829 4236422.919480448  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "558_1"
631096.2139024991 4236465.965779391  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "559_0"
648229.3396924527 4201793.2618079  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "560_0"
648042.0945841146 4201599.377172472  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "561_0"
647723.8863440289 4201568.264831236  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "561_1"
647469.9792322537 4201732.327952368  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "561_2"
646475.4809778115 4201690.279038115  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "561_3"
597912.6312819726 4215540.009304728  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "565_0"
597912.6312819726 4215540.009304728  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "566_0"
592434.7009135431 4213294.721300913  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "570_0"
591723.5130233101 4213839.196185748  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "570_1"
591013.9853944229 4214042.819844068  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "570_2"
590097.1608828605 4214301.361784798  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "571_0"
589099.7059368857 4214953.753904554  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "571_1"
588159.7876515206 4215151.995485564  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "571_2"
587333.2344210331 4219592.268165682  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "572_0"
585050.9027590858 4218980.703771464  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "572_1"
584245.8180855216 4218623.508769882  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "572_2"
586277.2663573823 4216988.988820302  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "573_0"
587270.0241211994 4217523.52520225  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "573_1"
588232.0405859168 4218057.753869937  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "573_2"
595026.5934640203 4214779.35433711  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "574_0"
593992.0590598079 4214184.641507439  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "574_1"
592975.7998466796 4213741.085326748  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "574_2"
591837.7790230004 4213128.655178311  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "574_3"
595042.9012020007 4214194.349763053  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "575_0"
594905.4010832546 4213461.407629166  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "575_1"
594309.7646466774 4212545.112558938  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "575_2"
593622.5972057834 4212407.619389435  0 0 "Arial" -11 0 0 0 0 0 0 0 0 0 0 0 0 "575_3"
